module udma_subsystem_tb;


	
endmodule