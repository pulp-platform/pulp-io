package pulp_io_pkg;
	
	
endpackage