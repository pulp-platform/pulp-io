`define HYPER_MACRO 1